module stop_cache

	(input do_replace,
	 input do_prop_write,
	 input mem_valid,

	 output stop_cache);


endmodule
